<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>16.488,5.54313,149.838,-66.2319</PageViewport>
<gate>
<ID>2</ID>
<type>AI_MUX_8x1</type>
<position>44.5,-24.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>5 </input>
<input>
<ID>IN_4</ID>4 </input>
<input>
<ID>IN_5</ID>3 </input>
<input>
<ID>IN_6</ID>2 </input>
<input>
<ID>IN_7</ID>1 </input>
<output>
<ID>OUT</ID>12 </output>
<input>
<ID>SEL_0</ID>11 </input>
<input>
<ID>SEL_1</ID>10 </input>
<input>
<ID>SEL_2</ID>9 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>23,-16.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>22.5,-19</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>22.5,-21.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>22.5,-24</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>22.5,-26.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>22.5,-29</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>22.5,-31.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>22,-34</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>42.5,-9.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>40.5,-12.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>39.5,-15.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>56.5,-24.5</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>BE_DECODER_3x8</type>
<position>42,-43</position>
<input>
<ID>ENABLE</ID>16 </input>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>13 </input>
<output>
<ID>OUT_0</ID>24 </output>
<output>
<ID>OUT_1</ID>23 </output>
<output>
<ID>OUT_2</ID>22 </output>
<output>
<ID>OUT_3</ID>21 </output>
<output>
<ID>OUT_4</ID>20 </output>
<output>
<ID>OUT_5</ID>19 </output>
<output>
<ID>OUT_6</ID>18 </output>
<output>
<ID>OUT_7</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>25,-43.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>25,-46.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>25,-49.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>27.5,-39</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>54.5,-39.5</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>GA_LED</type>
<position>54.5,-42</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>54.5,-44.5</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>GA_LED</type>
<position>54.5,-47</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>54.5,-49.5</position>
<input>
<ID>N_in0</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>54.5,-52</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>54.5,-54.5</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>54.5,-57</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>87,-30.5</position>
<output>
<ID>A_equal_B</ID>40 </output>
<output>
<ID>A_greater_B</ID>39 </output>
<output>
<ID>A_less_B</ID>41 </output>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<input>
<ID>IN_2</ID>26 </input>
<input>
<ID>IN_3</ID>25 </input>
<input>
<ID>IN_B_0</ID>32 </input>
<input>
<ID>IN_B_1</ID>31 </input>
<input>
<ID>IN_B_2</ID>30 </input>
<input>
<ID>IN_B_3</ID>29 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_TOGGLE</type>
<position>82.5,-18</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>85,-18</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>80,-18</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>77.5,-18</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>94,-18</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>96.5,-18</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>91.5,-18</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>89,-18</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>60</ID>
<type>GA_LED</type>
<position>72.5,-28.5</position>
<input>
<ID>N_in1</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>GA_LED</type>
<position>72.5,-31</position>
<input>
<ID>N_in1</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>72.5,-33.5</position>
<input>
<ID>N_in1</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-21,30.5,-16.5</points>
<intersection>-21 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-21,41.5,-21</points>
<connection>
<GID>2</GID>
<name>IN_7</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-16.5,30.5,-16.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-22,30.5,-19</points>
<intersection>-22 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-22,41.5,-22</points>
<connection>
<GID>2</GID>
<name>IN_6</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-19,30.5,-19</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-23,30.5,-21.5</points>
<intersection>-23 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-23,41.5,-23</points>
<connection>
<GID>2</GID>
<name>IN_5</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-21.5,30.5,-21.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-24,41.5,-24</points>
<connection>
<GID>2</GID>
<name>IN_4</name></connection>
<intersection>24.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>24.5,-24,24.5,-24</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-26.5,32,-25</points>
<intersection>-26.5 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-25,41.5,-25</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-26.5,32,-26.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-29,32,-26</points>
<intersection>-29 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-26,41.5,-26</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-29,32,-29</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-31.5,32,-27</points>
<intersection>-31.5 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-27,41.5,-27</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24.5,-31.5,32,-31.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-34,32,-28</points>
<intersection>-34 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-28,41.5,-28</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-34,32,-34</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-19,43.5,-15.5</points>
<connection>
<GID>2</GID>
<name>SEL_2</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-15.5,43.5,-15.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-19,44.5,-12.5</points>
<connection>
<GID>2</GID>
<name>SEL_1</name></connection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-12.5,44.5,-12.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-19,45.5,-9.5</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-9.5,45.5,-9.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,-24.5,55.5,-24.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>55.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>55.5,-24.5,55.5,-24.5</points>
<connection>
<GID>19</GID>
<name>N_in0</name></connection>
<intersection>-24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-44.5,34,-43.5</points>
<intersection>-44.5 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-44.5,39,-44.5</points>
<connection>
<GID>21</GID>
<name>IN_2</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-43.5,34,-43.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-46.5,33,-45.5</points>
<intersection>-46.5 2</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-45.5,39,-45.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-46.5,33,-46.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-49.5,32.5,-46.5</points>
<intersection>-49.5 2</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-46.5,39,-46.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-49.5,32.5,-49.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-39.5,39,-39.5</points>
<connection>
<GID>21</GID>
<name>ENABLE</name></connection>
<intersection>29.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29.5,-39.5,29.5,-39</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45,-39.5,53.5,-39.5</points>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<connection>
<GID>21</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-42,49,-40.5</points>
<intersection>-42 1</intersection>
<intersection>-40.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-42,53.5,-42</points>
<connection>
<GID>29</GID>
<name>N_in0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-40.5,49,-40.5</points>
<connection>
<GID>21</GID>
<name>OUT_6</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-44.5,49,-41.5</points>
<intersection>-44.5 1</intersection>
<intersection>-41.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-44.5,53.5,-44.5</points>
<connection>
<GID>30</GID>
<name>N_in0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-41.5,49,-41.5</points>
<connection>
<GID>21</GID>
<name>OUT_5</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-47,49,-42.5</points>
<intersection>-47 1</intersection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-47,53.5,-47</points>
<connection>
<GID>31</GID>
<name>N_in0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-42.5,49,-42.5</points>
<connection>
<GID>21</GID>
<name>OUT_4</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-49.5,49,-43.5</points>
<intersection>-49.5 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-49.5,53.5,-49.5</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-43.5,49,-43.5</points>
<connection>
<GID>21</GID>
<name>OUT_3</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-52,49,-44.5</points>
<intersection>-52 1</intersection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-52,53.5,-52</points>
<connection>
<GID>33</GID>
<name>N_in0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-44.5,49,-44.5</points>
<connection>
<GID>21</GID>
<name>OUT_2</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-54.5,49,-45.5</points>
<intersection>-54.5 1</intersection>
<intersection>-45.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-54.5,53.5,-54.5</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-45.5,49,-45.5</points>
<connection>
<GID>21</GID>
<name>OUT_1</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-57,49,-46.5</points>
<intersection>-57 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-57,53.5,-57</points>
<connection>
<GID>35</GID>
<name>N_in0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45,-46.5,49,-46.5</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-26.5,82,-23</points>
<connection>
<GID>39</GID>
<name>IN_3</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>77.5,-23,77.5,-20</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-23,82,-23</points>
<intersection>77.5 1</intersection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-26.5,83,-23</points>
<connection>
<GID>39</GID>
<name>IN_2</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>80,-23,80,-20</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>80,-23,83,-23</points>
<intersection>80 1</intersection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-26.5,84,-23</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>82.5,-23,82.5,-20</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-23,84,-23</points>
<intersection>82.5 1</intersection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-26.5,85,-20</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>-26.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>85,-26.5,85,-26.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-26.5,89,-20</points>
<connection>
<GID>39</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-26.5,90,-23</points>
<connection>
<GID>39</GID>
<name>IN_B_2</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>91.5,-23,91.5,-20</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>90,-23,91.5,-23</points>
<intersection>90 0</intersection>
<intersection>91.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-26.5,91,-23</points>
<connection>
<GID>39</GID>
<name>IN_B_1</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>94,-23,94,-20</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91,-23,94,-23</points>
<intersection>91 0</intersection>
<intersection>94 1</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-26.5,92,-23</points>
<connection>
<GID>39</GID>
<name>IN_B_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>96.5,-23,96.5,-20</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>92,-23,96.5,-23</points>
<intersection>92 0</intersection>
<intersection>96.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-28.5,79,-28.5</points>
<connection>
<GID>60</GID>
<name>N_in1</name></connection>
<connection>
<GID>39</GID>
<name>A_greater_B</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-31,76,-30.5</points>
<intersection>-31 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-31,76,-31</points>
<connection>
<GID>61</GID>
<name>N_in1</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76,-30.5,79,-30.5</points>
<connection>
<GID>39</GID>
<name>A_equal_B</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-33.5,76,-32.5</points>
<intersection>-33.5 1</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-33.5,76,-33.5</points>
<connection>
<GID>62</GID>
<name>N_in1</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76,-32.5,79,-32.5</points>
<connection>
<GID>39</GID>
<name>A_less_B</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 9></circuit>