<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-57.762,5.54313,75.588,-66.2319</PageViewport>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>40.5,-18.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_OR2</type>
<position>52.5,-13.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_INVERTER</type>
<position>40.5,-10</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>28.5,-10.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>29,-17.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>29,-20.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>71,-13.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_INVERTER</type>
<position>62.5,-13.5</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_INVERTER</type>
<position>40.5,-43.5</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>40.5,-36</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>40.5,-30.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>27.5,-31</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>27.5,-34.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>28,-37.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AE_OR2</type>
<position>54,-39</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_OR2</type>
<position>63.5,-34.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>-38.5,-9</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>69,-34.5</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_INVERTER</type>
<position>-7.5,-17</position>
<input>
<ID>IN_0</ID>19 </input>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_INVERTER</type>
<position>-7.5,-21</position>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_TOGGLE</type>
<position>-38.5,-14</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>-38.5,-18.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_AND2</type>
<position>-29.5,-15.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>-26.5,-23.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>AE_OR2</type>
<position>-21,-10.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>AE_OR2</type>
<position>-19,-21</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_AND2</type>
<position>4,-19</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AE_OR2</type>
<position>-66,-6</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>GA_LED</type>
<position>10.5,-19</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-10.5,37.5,-10.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>37.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,-10.5,37.5,-10</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-17.5,37.5,-17.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>37.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,-17.5,37.5,-17.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-20.5,34,-19.5</points>
<intersection>-20.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-19.5,37.5,-19.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-20.5,34,-20.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-18.5,46.5,-14.5</points>
<intersection>-18.5 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-14.5,49.5,-14.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-18.5,46.5,-18.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-12.5,46.5,-10</points>
<intersection>-12.5 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-12.5,49.5,-12.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-10,46.5,-10</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55.5,-13.5,59.5,-13.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,-13.5,70,-13.5</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-31,33.5,-29.5</points>
<intersection>-31 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-29.5,37.5,-29.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-31,33.5,-31</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-34.5,33.5,-31.5</points>
<intersection>-34.5 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-31.5,37.5,-31.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>33.5 0</intersection>
<intersection>37.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-34.5,33.5,-34.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,-35,37.5,-31.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-31.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-37.5,33.5,-37</points>
<intersection>-37.5 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-37,37.5,-37</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>33.5 0</intersection>
<intersection>37.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-37.5,33.5,-37.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,-43.5,37.5,-37</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-37 1</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-33.5,52,-30.5</points>
<intersection>-33.5 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-33.5,60.5,-33.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-30.5,52,-30.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-38,47,-36</points>
<intersection>-38 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-38,51,-38</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-36,47,-36</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-43.5,47,-40</points>
<intersection>-43.5 2</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-40,51,-40</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-43.5,47,-43.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-39,58.5,-35.5</points>
<intersection>-39 2</intersection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-35.5,60.5,-35.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-39,58.5,-39</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,-34.5,68,-34.5</points>
<connection>
<GID>35</GID>
<name>N_in0</name></connection>
<connection>
<GID>31</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-24.5,-30,-9</points>
<intersection>-24.5 3</intersection>
<intersection>-9.5 1</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-9.5,-24,-9.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-36.5,-9,-30,-9</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-30,-24.5,-29.5,-24.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-17,-14,-10.5</points>
<intersection>-17 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-17,-10.5,-17</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-18,-10.5,-14,-10.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,-15.5,-25,-11.5</points>
<intersection>-15.5 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,-11.5,-24,-11.5</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-26.5,-15.5,-25,-15.5</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36.5,-14,-22,-14</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 4</intersection>
<intersection>-22 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-22,-20,-22,-14</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-32.5,-14.5,-32.5,-14</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34.5,-22.5,-34.5,-16.5</points>
<intersection>-22.5 3</intersection>
<intersection>-18.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-16.5,-32.5,-16.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>-34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-36.5,-18.5,-34.5,-18.5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>-34.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-34.5,-22.5,-29.5,-22.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>-34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22.5,-23.5,-22.5,-22</points>
<intersection>-23.5 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22.5,-22,-22,-22</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>-22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-23.5,-23.5,-22.5,-23.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>-22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16,-21,-10.5,-21</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<connection>
<GID>51</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-21,-1.5,-20</points>
<intersection>-21 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,-20,1,-20</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4.5,-21,-1.5,-21</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-18,-1.5,-17</points>
<intersection>-18 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,-18,1,-18</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4.5,-17,-1.5,-17</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-19,9.5,-19</points>
<connection>
<GID>57</GID>
<name>N_in0</name></connection>
<connection>
<GID>53</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-95.7</PageViewport></page 9></circuit>